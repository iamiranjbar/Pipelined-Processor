module adder(input[11:0] a,b,output logic[11:0] out);
  assign out=a+b;
endmodule
