module CU(input [4:0] func,input Z,C,rst,output logic ld_pc,push,pop,reg_write_en,sel1_ALU_in,sel2_ALU_in,ldzero,ldcarry,sel_second_load,mem_write_en,mem_read,sel_data_RF_write, output logic[1:0] instSel);
  always @(*)  
  begin 
  if(rst)begin
    ld_pc=1'b0;
    instSel=1'b0;
    push=1'b0;
    pop=1'b0;
    reg_write_en=1'b0;
    sel1_ALU_in=1'b0;
    sel2_ALU_in=1'b0;
    ldzero=1'b0;
    ldcarry=1'b0;
    sel_second_load=1'b0;
    mem_write_en=1'b0;
    mem_read=1'b0;
    sel_data_RF_write=1'b0;
  end
  else begin
    case(func)
      5'b00000:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b0;
        sel2_ALU_in=1'b0;
        ldzero=1'b1;
        ldcarry=1'b1;
        sel_data_RF_write=1'b1;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b00001:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b0;
        sel2_ALU_in=1'b0;
        ldzero=1'b1;
        ldcarry=1'b1;
        sel_data_RF_write=1'b1;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b00010:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b0;
        sel2_ALU_in=1'b0;
        ldzero=1'b1;
        ldcarry=1'b1;
        sel_data_RF_write=1'b1;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b00011:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b0;
        sel2_ALU_in=1'b0;
        ldzero=1'b1;
        ldcarry=1'b1;
        sel_data_RF_write=1'b1;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b00100:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b0;
        sel2_ALU_in=1'b0;
        ldzero=1'b1;
        ldcarry=1'b1;
        sel_data_RF_write=1'b1;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b00101:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b0;
        sel2_ALU_in=1'b0;
        ldzero=1'b1;
        ldcarry=1'b1;
        sel_data_RF_write=1'b1;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b00110:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b0;
        sel2_ALU_in=1'b0;
        ldzero=1'b1;
        ldcarry=1'b1;
        sel_data_RF_write=1'b1;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b00111:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b0;
        sel2_ALU_in=1'b0;
        ldzero=1'b1;
        ldcarry=1'b1;
        sel_data_RF_write=1'b1;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b01000:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b1;
        sel2_ALU_in=1'b0;
        ldzero=1'b1;
        ldcarry=1'b1;
        sel_data_RF_write=1'b1;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b01001:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b1;
        sel2_ALU_in=1'b0;
        ldzero=1'b1;
        ldcarry=1'b1;
        sel_data_RF_write=1'b1;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b01010:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b1;
        sel2_ALU_in=1'b0;
        ldzero=1'b1;
        ldcarry=1'b1;
        sel_data_RF_write=1'b1;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b01011:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b1;
        sel2_ALU_in=1'b0;
        ldzero=1'b1;
        ldcarry=1'b1;
        sel_data_RF_write=1'b1;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b01100:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b1;
        sel2_ALU_in=1'b0;
        ldzero=1'b1;
        ldcarry=1'b1;
        sel_data_RF_write=1'b1;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b01101:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b1;
        sel2_ALU_in=1'b0;
        ldzero=1'b1;
        ldcarry=1'b1;
        sel_data_RF_write=1'b1;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b01110:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b1;
        sel2_ALU_in=1'b0;
        ldzero=1'b1;
        ldcarry=1'b1;
        sel_data_RF_write=1'b1;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b01111:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b1;
        sel2_ALU_in=1'b0;
        ldzero=1'b1;
        ldcarry=1'b1;
        sel_data_RF_write=1'b1;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b11000:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b0;
        sel2_ALU_in=1'b1;
        ldzero=1'b1;
        ldcarry=1'b1;
        sel_data_RF_write=1'b1;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b11001:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b0;
        sel2_ALU_in=1'b1;
        ldzero=1'b1;
        ldcarry=1'b1;
        sel_data_RF_write=1'b1;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b11010:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b0;
        sel2_ALU_in=1'b1;
        ldzero=1'b1;
        ldcarry=1'b1;
        sel_data_RF_write=1'b1;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b11011:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b0;
        sel2_ALU_in=1'b1;
        ldzero=1'b1;
        ldcarry=1'b1;
        sel_data_RF_write=1'b1;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b10000:begin
        instSel=1'b1;
        sel_second_load=1'b1;
        sel1_ALU_in=1'b1;
        sel2_ALU_in=1'b0;
        ldzero=1'b0;
        ldcarry=1'b0;
        sel_data_RF_write=1'b0;
        reg_write_en=1'b1;
        mem_write_en=1'b0;
        mem_read=1'b1;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b10001:begin
        instSel=1'b1;
        sel_second_load=1'b0;
        sel1_ALU_in=1'b1;
        sel2_ALU_in=1'b0;
        ldzero=1'b0;
        ldcarry=1'b0;
        sel_data_RF_write=1'b0;
        reg_write_en=1'b0;
        mem_write_en=1'b1;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b10100:begin
        instSel=(Z)?1'b0:1'b1;
        sel_second_load=1'b0;
        sel1_ALU_in=1'b0;
        sel2_ALU_in=1'b0;
        ldzero=1'b0;
        ldcarry=1'b0;
        sel_data_RF_write=1'b0;
        reg_write_en=1'b0;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b10101:begin
        instSel=(~Z)?1'b0:1'b1;
        sel_second_load=1'b0;
        sel1_ALU_in=1'b0;
        sel2_ALU_in=1'b0;
        ldzero=1'b0;
        ldcarry=1'b0;
        sel_data_RF_write=1'b0;
        reg_write_en=1'b0;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b10110:begin
        instSel=(C)?1'b0:1'b1;
        sel_second_load=1'b0;
        sel1_ALU_in=1'b0;
        sel2_ALU_in=1'b0;
        ldzero=1'b0;
        ldcarry=1'b0;
        sel_data_RF_write=1'b0;
        reg_write_en=1'b0;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b10111:begin
        instSel=(~C)?1'b0:1'b1;
        sel_second_load=1'b0;
        sel1_ALU_in=1'b0;
        sel2_ALU_in=1'b0;
        ldzero=1'b0;
        ldcarry=1'b0;
        sel_data_RF_write=1'b0;
        reg_write_en=1'b0;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b11100:begin
        instSel=1'b1;
        sel_second_load=1'b0;
        sel1_ALU_in=1'b0;
        sel2_ALU_in=1'b0;
        ldzero=1'b0;
        ldcarry=1'b0;
        sel_data_RF_write=1'b0;
        reg_write_en=1'b0;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b11101:begin
        instSel=1'b1;
        sel_second_load=1'b0;
        sel1_ALU_in=1'b0;
        sel2_ALU_in=1'b0;
        ldzero=1'b0;
        ldcarry=1'b0;
        sel_data_RF_write=1'b0;
        reg_write_en=1'b0;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b1;
        pop=1'b0;
        ld_pc=1'b1;
      end
      5'b11110:begin
        instSel=1'b1;
        sel_second_load=1'b0;
        sel1_ALU_in=1'b0;
        sel2_ALU_in=1'b0;
        ldzero=1'b0;
        ldcarry=1'b0;
        sel_data_RF_write=1'b0;
        reg_write_en=1'b0;
        mem_write_en=1'b0;
        mem_read=1'b0;
        push=1'b0;
        pop=1'b1;
        ld_pc=1'b1;
      end
    endcase
  end
  end
endmodule
