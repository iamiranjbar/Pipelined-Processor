module flushMux();

endmodule