module flushDetection(input ID_EX_memRead, input [2:0] Rs, Rt, ID_EX_Rt, output flushMuxSel, PCWr, IF_ID_Wr);
	
endmodule